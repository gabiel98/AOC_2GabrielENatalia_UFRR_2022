-- Somador do PC
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SomadorPC IS
PORT(
	   SomaIn 					: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		Soma2						: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		SomaOut 					: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));

END SomadorPC;

ARCHITECTURE behavior OF SomadorPC IS
BEGIN
	SomaOut <= SomaIn + Soma2;
	
END behavior;